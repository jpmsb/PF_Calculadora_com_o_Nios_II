-- system.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		clk_clk                                : in    std_logic                     := '0';             --                             clk.clk
		entrada_pio_external_connection_export : in    std_logic_vector(18 downto 0) := (others => '0'); -- entrada_pio_external_connection.export
		lcd_16x2_external_interface_DATA       : inout std_logic_vector(7 downto 0)  := (others => '0'); --     lcd_16x2_external_interface.DATA
		lcd_16x2_external_interface_ON         : out   std_logic;                                        --                                .ON
		lcd_16x2_external_interface_BLON       : out   std_logic;                                        --                                .BLON
		lcd_16x2_external_interface_EN         : out   std_logic;                                        --                                .EN
		lcd_16x2_external_interface_RS         : out   std_logic;                                        --                                .RS
		lcd_16x2_external_interface_RW         : out   std_logic;                                        --                                .RW
		led_pio_external_connection_export     : out   std_logic_vector(15 downto 0);                    --     led_pio_external_connection.export
		reset_reset_n                          : in    std_logic                     := '0'              --                           reset.reset_n
	);
end entity system;

architecture rtl of system is
	component system_entrada_pio is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(18 downto 0) := (others => 'X')  -- export
		);
	end component system_entrada_pio;

	component system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_jtag_uart;

	component system_lcd_16x2 is
		port (
			clk         : in    std_logic                    := 'X';             -- clk
			reset       : in    std_logic                    := 'X';             -- reset
			address     : in    std_logic                    := 'X';             -- address
			chipselect  : in    std_logic                    := 'X';             -- chipselect
			read        : in    std_logic                    := 'X';             -- read
			write       : in    std_logic                    := 'X';             -- write
			writedata   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(7 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                       -- waitrequest
			LCD_DATA    : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_ON      : out   std_logic;                                       -- export
			LCD_BLON    : out   std_logic;                                       -- export
			LCD_EN      : out   std_logic;                                       -- export
			LCD_RS      : out   std_logic;                                       -- export
			LCD_RW      : out   std_logic                                        -- export
		);
	end component system_lcd_16x2;

	component system_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component system_led_pio;

	component system_nios2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_nios2_0;

	component system_onchip_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component system_onchip_mem;

	component system_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component system_sys_clk_timer;

	component system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component system_sysid;

	component system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			nios2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_0_data_master_address               : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			nios2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_0_data_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			nios2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_0_instruction_master_address        : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			nios2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_0_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			entrada_pio_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			entrada_pio_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_address       : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write         : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read          : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect    : out std_logic;                                        -- chipselect
			lcd_16x2_avalon_lcd_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			lcd_16x2_avalon_lcd_slave_write           : out std_logic;                                        -- write
			lcd_16x2_avalon_lcd_slave_read            : out std_logic;                                        -- read
			lcd_16x2_avalon_lcd_slave_readdata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			lcd_16x2_avalon_lcd_slave_writedata       : out std_logic_vector(7 downto 0);                     -- writedata
			lcd_16x2_avalon_lcd_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			lcd_16x2_avalon_lcd_slave_chipselect      : out std_logic;                                        -- chipselect
			led_pio_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                          : out std_logic;                                        -- write
			led_pio_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                     : out std_logic;                                        -- chipselect
			nios2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			onchip_mem_s1_address                     : out std_logic_vector(13 downto 0);                    -- address
			onchip_mem_s1_write                       : out std_logic;                                        -- write
			onchip_mem_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_mem_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_mem_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_mem_s1_chipselect                  : out std_logic;                                        -- chipselect
			onchip_mem_s1_clken                       : out std_logic;                                        -- clken
			sys_clk_timer_s1_address                  : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                    : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect               : out std_logic;                                        -- chipselect
			sysid_control_slave_address               : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_0_data_master_readdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_0_data_master_readdata -> nios2_0:d_readdata
	signal nios2_0_data_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:nios2_0_data_master_waitrequest -> nios2_0:d_waitrequest
	signal nios2_0_data_master_debugaccess                               : std_logic;                     -- nios2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_0_data_master_debugaccess
	signal nios2_0_data_master_address                                   : std_logic_vector(17 downto 0); -- nios2_0:d_address -> mm_interconnect_0:nios2_0_data_master_address
	signal nios2_0_data_master_byteenable                                : std_logic_vector(3 downto 0);  -- nios2_0:d_byteenable -> mm_interconnect_0:nios2_0_data_master_byteenable
	signal nios2_0_data_master_read                                      : std_logic;                     -- nios2_0:d_read -> mm_interconnect_0:nios2_0_data_master_read
	signal nios2_0_data_master_readdatavalid                             : std_logic;                     -- mm_interconnect_0:nios2_0_data_master_readdatavalid -> nios2_0:d_readdatavalid
	signal nios2_0_data_master_write                                     : std_logic;                     -- nios2_0:d_write -> mm_interconnect_0:nios2_0_data_master_write
	signal nios2_0_data_master_writedata                                 : std_logic_vector(31 downto 0); -- nios2_0:d_writedata -> mm_interconnect_0:nios2_0_data_master_writedata
	signal nios2_0_instruction_master_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_0_instruction_master_readdata -> nios2_0:i_readdata
	signal nios2_0_instruction_master_waitrequest                        : std_logic;                     -- mm_interconnect_0:nios2_0_instruction_master_waitrequest -> nios2_0:i_waitrequest
	signal nios2_0_instruction_master_address                            : std_logic_vector(17 downto 0); -- nios2_0:i_address -> mm_interconnect_0:nios2_0_instruction_master_address
	signal nios2_0_instruction_master_read                               : std_logic;                     -- nios2_0:i_read -> mm_interconnect_0:nios2_0_instruction_master_read
	signal nios2_0_instruction_master_readdatavalid                      : std_logic;                     -- mm_interconnect_0:nios2_0_instruction_master_readdatavalid -> nios2_0:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_lcd_16x2_avalon_lcd_slave_chipselect        : std_logic;                     -- mm_interconnect_0:lcd_16x2_avalon_lcd_slave_chipselect -> lcd_16x2:chipselect
	signal mm_interconnect_0_lcd_16x2_avalon_lcd_slave_readdata          : std_logic_vector(7 downto 0);  -- lcd_16x2:readdata -> mm_interconnect_0:lcd_16x2_avalon_lcd_slave_readdata
	signal mm_interconnect_0_lcd_16x2_avalon_lcd_slave_waitrequest       : std_logic;                     -- lcd_16x2:waitrequest -> mm_interconnect_0:lcd_16x2_avalon_lcd_slave_waitrequest
	signal mm_interconnect_0_lcd_16x2_avalon_lcd_slave_address           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:lcd_16x2_avalon_lcd_slave_address -> lcd_16x2:address
	signal mm_interconnect_0_lcd_16x2_avalon_lcd_slave_read              : std_logic;                     -- mm_interconnect_0:lcd_16x2_avalon_lcd_slave_read -> lcd_16x2:read
	signal mm_interconnect_0_lcd_16x2_avalon_lcd_slave_write             : std_logic;                     -- mm_interconnect_0:lcd_16x2_avalon_lcd_slave_write -> lcd_16x2:write
	signal mm_interconnect_0_lcd_16x2_avalon_lcd_slave_writedata         : std_logic_vector(7 downto 0);  -- mm_interconnect_0:lcd_16x2_avalon_lcd_slave_writedata -> lcd_16x2:writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_nios2_0_debug_mem_slave_readdata            : std_logic_vector(31 downto 0); -- nios2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest         : std_logic;                     -- nios2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess         : std_logic;                     -- mm_interconnect_0:nios2_0_debug_mem_slave_debugaccess -> nios2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_0_debug_mem_slave_address             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_0_debug_mem_slave_address -> nios2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_0_debug_mem_slave_read                : std_logic;                     -- mm_interconnect_0:nios2_0_debug_mem_slave_read -> nios2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_0_debug_mem_slave_byteenable          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_0_debug_mem_slave_byteenable -> nios2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_0_debug_mem_slave_write               : std_logic;                     -- mm_interconnect_0:nios2_0_debug_mem_slave_write -> nios2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_0_debug_mem_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_0_debug_mem_slave_writedata -> nios2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_led_pio_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_0_led_pio_s1_readdata                         : std_logic_vector(31 downto 0); -- led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	signal mm_interconnect_0_led_pio_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_0_led_pio_s1_write                            : std_logic;                     -- mm_interconnect_0:led_pio_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	signal mm_interconnect_0_onchip_mem_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	signal mm_interconnect_0_onchip_mem_s1_readdata                      : std_logic_vector(31 downto 0); -- onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	signal mm_interconnect_0_onchip_mem_s1_address                       : std_logic_vector(13 downto 0); -- mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	signal mm_interconnect_0_onchip_mem_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	signal mm_interconnect_0_onchip_mem_s1_write                         : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	signal mm_interconnect_0_onchip_mem_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	signal mm_interconnect_0_onchip_mem_s1_clken                         : std_logic;                     -- mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	signal mm_interconnect_0_sys_clk_timer_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_0_sys_clk_timer_s1_readdata                   : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	signal mm_interconnect_0_sys_clk_timer_s1_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_0_sys_clk_timer_s1_write                      : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_write -> mm_interconnect_0_sys_clk_timer_s1_write:in
	signal mm_interconnect_0_sys_clk_timer_s1_writedata                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_0_entrada_pio_s1_readdata                     : std_logic_vector(31 downto 0); -- entrada_pio:readdata -> mm_interconnect_0:entrada_pio_s1_readdata
	signal mm_interconnect_0_entrada_pio_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:entrada_pio_s1_address -> entrada_pio:address
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver1_irq
	signal nios2_0_irq_irq                                               : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_0:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, lcd_16x2:reset, mm_interconnect_0:nios2_0_reset_reset_bridge_in_reset_reset, onchip_mem:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [nios2_0:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_led_pio_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_led_pio_s1_write:inv -> led_pio:write_n
	signal mm_interconnect_0_sys_clk_timer_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [entrada_pio:reset_n, jtag_uart:rst_n, led_pio:reset_n, nios2_0:reset_n, sys_clk_timer:reset_n, sysid:reset_n]

begin

	entrada_pio : component system_entrada_pio
		port map (
			clk      => clk_clk,                                   --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => mm_interconnect_0_entrada_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_entrada_pio_s1_readdata, --                    .readdata
			in_port  => entrada_pio_external_connection_export     -- external_connection.export
		);

	jtag_uart : component system_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	lcd_16x2 : component system_lcd_16x2
		port map (
			clk         => clk_clk,                                                 --                clk.clk
			reset       => rst_controller_reset_out_reset,                          --              reset.reset
			address     => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_address(0),  --   avalon_lcd_slave.address
			chipselect  => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_chipselect,  --                   .chipselect
			read        => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_read,        --                   .read
			write       => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_write,       --                   .write
			writedata   => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_waitrequest, --                   .waitrequest
			LCD_DATA    => lcd_16x2_external_interface_DATA,                        -- external_interface.export
			LCD_ON      => lcd_16x2_external_interface_ON,                          --                   .export
			LCD_BLON    => lcd_16x2_external_interface_BLON,                        --                   .export
			LCD_EN      => lcd_16x2_external_interface_EN,                          --                   .export
			LCD_RS      => lcd_16x2_external_interface_RS,                          --                   .export
			LCD_RW      => lcd_16x2_external_interface_RW                           --                   .export
		);

	led_pio : component system_led_pio
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	nios2_0 : component system_nios2_0
		port map (
			clk                                 => clk_clk,                                               --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,              --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                           => nios2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                  --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                   -- custom_instruction_master.readra
		);

	onchip_mem : component system_onchip_mem
		port map (
			clk        => clk_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	sys_clk_timer : component system_sys_clk_timer
		port map (
			clk        => clk_clk,                                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                            --   irq.irq
		);

	sysid : component system_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                                   --                           clk_0_clk.clk
			nios2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- nios2_0_reset_reset_bridge_in_reset.reset
			nios2_0_data_master_address               => nios2_0_data_master_address,                               --                 nios2_0_data_master.address
			nios2_0_data_master_waitrequest           => nios2_0_data_master_waitrequest,                           --                                    .waitrequest
			nios2_0_data_master_byteenable            => nios2_0_data_master_byteenable,                            --                                    .byteenable
			nios2_0_data_master_read                  => nios2_0_data_master_read,                                  --                                    .read
			nios2_0_data_master_readdata              => nios2_0_data_master_readdata,                              --                                    .readdata
			nios2_0_data_master_readdatavalid         => nios2_0_data_master_readdatavalid,                         --                                    .readdatavalid
			nios2_0_data_master_write                 => nios2_0_data_master_write,                                 --                                    .write
			nios2_0_data_master_writedata             => nios2_0_data_master_writedata,                             --                                    .writedata
			nios2_0_data_master_debugaccess           => nios2_0_data_master_debugaccess,                           --                                    .debugaccess
			nios2_0_instruction_master_address        => nios2_0_instruction_master_address,                        --          nios2_0_instruction_master.address
			nios2_0_instruction_master_waitrequest    => nios2_0_instruction_master_waitrequest,                    --                                    .waitrequest
			nios2_0_instruction_master_read           => nios2_0_instruction_master_read,                           --                                    .read
			nios2_0_instruction_master_readdata       => nios2_0_instruction_master_readdata,                       --                                    .readdata
			nios2_0_instruction_master_readdatavalid  => nios2_0_instruction_master_readdatavalid,                  --                                    .readdatavalid
			entrada_pio_s1_address                    => mm_interconnect_0_entrada_pio_s1_address,                  --                      entrada_pio_s1.address
			entrada_pio_s1_readdata                   => mm_interconnect_0_entrada_pio_s1_readdata,                 --                                    .readdata
			jtag_uart_avalon_jtag_slave_address       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --         jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                    .write
			jtag_uart_avalon_jtag_slave_read          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                    .read
			jtag_uart_avalon_jtag_slave_readdata      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                    .readdata
			jtag_uart_avalon_jtag_slave_writedata     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                    .writedata
			jtag_uart_avalon_jtag_slave_waitrequest   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                    .chipselect
			lcd_16x2_avalon_lcd_slave_address         => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_address,       --           lcd_16x2_avalon_lcd_slave.address
			lcd_16x2_avalon_lcd_slave_write           => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_write,         --                                    .write
			lcd_16x2_avalon_lcd_slave_read            => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_read,          --                                    .read
			lcd_16x2_avalon_lcd_slave_readdata        => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_readdata,      --                                    .readdata
			lcd_16x2_avalon_lcd_slave_writedata       => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_writedata,     --                                    .writedata
			lcd_16x2_avalon_lcd_slave_waitrequest     => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_waitrequest,   --                                    .waitrequest
			lcd_16x2_avalon_lcd_slave_chipselect      => mm_interconnect_0_lcd_16x2_avalon_lcd_slave_chipselect,    --                                    .chipselect
			led_pio_s1_address                        => mm_interconnect_0_led_pio_s1_address,                      --                          led_pio_s1.address
			led_pio_s1_write                          => mm_interconnect_0_led_pio_s1_write,                        --                                    .write
			led_pio_s1_readdata                       => mm_interconnect_0_led_pio_s1_readdata,                     --                                    .readdata
			led_pio_s1_writedata                      => mm_interconnect_0_led_pio_s1_writedata,                    --                                    .writedata
			led_pio_s1_chipselect                     => mm_interconnect_0_led_pio_s1_chipselect,                   --                                    .chipselect
			nios2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_0_debug_mem_slave_address,         --             nios2_0_debug_mem_slave.address
			nios2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_0_debug_mem_slave_write,           --                                    .write
			nios2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_0_debug_mem_slave_read,            --                                    .read
			nios2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_0_debug_mem_slave_readdata,        --                                    .readdata
			nios2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_0_debug_mem_slave_writedata,       --                                    .writedata
			nios2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_0_debug_mem_slave_byteenable,      --                                    .byteenable
			nios2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_0_debug_mem_slave_waitrequest,     --                                    .waitrequest
			nios2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_0_debug_mem_slave_debugaccess,     --                                    .debugaccess
			onchip_mem_s1_address                     => mm_interconnect_0_onchip_mem_s1_address,                   --                       onchip_mem_s1.address
			onchip_mem_s1_write                       => mm_interconnect_0_onchip_mem_s1_write,                     --                                    .write
			onchip_mem_s1_readdata                    => mm_interconnect_0_onchip_mem_s1_readdata,                  --                                    .readdata
			onchip_mem_s1_writedata                   => mm_interconnect_0_onchip_mem_s1_writedata,                 --                                    .writedata
			onchip_mem_s1_byteenable                  => mm_interconnect_0_onchip_mem_s1_byteenable,                --                                    .byteenable
			onchip_mem_s1_chipselect                  => mm_interconnect_0_onchip_mem_s1_chipselect,                --                                    .chipselect
			onchip_mem_s1_clken                       => mm_interconnect_0_onchip_mem_s1_clken,                     --                                    .clken
			sys_clk_timer_s1_address                  => mm_interconnect_0_sys_clk_timer_s1_address,                --                    sys_clk_timer_s1.address
			sys_clk_timer_s1_write                    => mm_interconnect_0_sys_clk_timer_s1_write,                  --                                    .write
			sys_clk_timer_s1_readdata                 => mm_interconnect_0_sys_clk_timer_s1_readdata,               --                                    .readdata
			sys_clk_timer_s1_writedata                => mm_interconnect_0_sys_clk_timer_s1_writedata,              --                                    .writedata
			sys_clk_timer_s1_chipselect               => mm_interconnect_0_sys_clk_timer_s1_chipselect,             --                                    .chipselect
			sysid_control_slave_address               => mm_interconnect_0_sysid_control_slave_address,             --                 sysid_control_slave.address
			sysid_control_slave_readdata              => mm_interconnect_0_sysid_control_slave_readdata             --                                    .readdata
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_0_irq_irq                 --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	mm_interconnect_0_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_timer_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of system
